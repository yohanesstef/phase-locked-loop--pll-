magic
tech sky130A
timestamp 1717263486
<< metal1 >>
rect -115 1432 694 1472
rect -115 -698 -15 1432
rect 145 1414 795 1417
rect 144 1377 795 1414
rect 144 1051 244 1377
rect 350 1111 387 1156
rect 350 1081 353 1111
rect 384 1081 387 1111
rect 350 1078 387 1081
rect 1543 1063 1578 1100
rect 1543 1060 1579 1063
rect 144 951 245 1051
rect 1543 1030 1546 1060
rect 1576 1030 1579 1060
rect 1543 1027 1579 1030
rect 1956 1060 2056 1063
rect 1956 1030 1960 1060
rect 2052 1030 2056 1060
rect 145 13 245 951
rect 145 -87 460 13
rect 355 -498 460 -492
rect 355 -530 360 -498
rect 450 -530 460 -498
rect 355 -600 460 -530
rect 946 -698 1046 -548
rect -115 -798 1046 -698
rect 1108 -698 1208 -549
rect 1956 -698 2056 1030
rect 1108 -798 2056 -698
<< via1 >>
rect 353 1081 384 1111
rect 1546 1030 1576 1060
rect 1960 1030 2052 1060
rect 360 -530 450 -498
<< metal2 >>
rect 350 1111 387 1114
rect 350 1081 353 1111
rect 384 1081 387 1111
rect 350 1012 387 1081
rect 1543 1060 2056 1063
rect 1543 1030 1546 1060
rect 1576 1030 1960 1060
rect 2052 1030 2056 1060
rect 1543 1027 2056 1030
rect 350 -498 459 1012
rect 350 -530 360 -498
rect 450 -530 459 -498
rect 350 -599 459 -530
use pfd_ver4  pfd_ver4_0
timestamp 1717247908
transform 1 0 175 0 1 -251
box 185 -398 1676 264
use vco  vco_0
timestamp 1717262165
transform 1 0 258 0 1 817
box -300 -855 1950 1775
<< end >>
