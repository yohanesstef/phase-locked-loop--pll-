magic
tech sky130A
timestamp 1717262165
<< isosubstrate >>
rect 190 315 210 335
rect 400 325 405 345
rect 420 340 470 345
rect 420 325 490 340
rect 470 320 490 325
rect 715 315 770 355
rect 960 325 965 345
rect 980 340 1030 345
rect 980 325 1050 340
rect 1030 320 1050 325
rect 1275 315 1330 355
rect 1520 325 1525 345
rect 1540 340 1590 345
rect 1540 325 1610 340
rect 1590 320 1610 325
<< nwell >>
rect 60 460 210 625
rect 340 460 490 625
rect 620 460 770 625
rect 900 460 1050 625
rect 1180 460 1330 625
rect 1460 460 1610 625
<< nmos >>
rect 125 380 145 425
rect 405 380 425 425
rect 685 380 705 425
rect 965 380 985 425
rect 1245 380 1265 425
rect 1525 380 1545 425
<< pmos >>
rect 125 490 145 535
rect 405 490 425 535
rect 685 490 705 535
rect 965 490 985 535
rect 1245 490 1265 535
rect 1525 490 1545 535
<< ndiff >>
rect 80 420 125 425
rect 80 385 90 420
rect 110 385 125 420
rect 80 380 125 385
rect 145 420 190 425
rect 145 385 160 420
rect 180 385 190 420
rect 145 380 190 385
rect 360 420 405 425
rect 360 385 370 420
rect 390 385 405 420
rect 360 380 405 385
rect 425 420 470 425
rect 425 385 440 420
rect 460 385 470 420
rect 425 380 470 385
rect 640 420 685 425
rect 640 385 650 420
rect 670 385 685 420
rect 640 380 685 385
rect 705 420 750 425
rect 705 385 720 420
rect 740 385 750 420
rect 705 380 750 385
rect 920 420 965 425
rect 920 385 930 420
rect 950 385 965 420
rect 920 380 965 385
rect 985 420 1030 425
rect 985 385 1000 420
rect 1020 385 1030 420
rect 985 380 1030 385
rect 1200 420 1245 425
rect 1200 385 1210 420
rect 1230 385 1245 420
rect 1200 380 1245 385
rect 1265 420 1310 425
rect 1265 385 1280 420
rect 1300 385 1310 420
rect 1265 380 1310 385
rect 1480 420 1525 425
rect 1480 385 1490 420
rect 1510 385 1525 420
rect 1480 380 1525 385
rect 1545 420 1590 425
rect 1545 385 1560 420
rect 1580 385 1590 420
rect 1545 380 1590 385
<< pdiff >>
rect 80 530 125 535
rect 80 495 90 530
rect 110 495 125 530
rect 80 490 125 495
rect 145 530 190 535
rect 145 495 160 530
rect 180 495 190 530
rect 145 490 190 495
rect 360 530 405 535
rect 360 495 370 530
rect 390 495 405 530
rect 360 490 405 495
rect 425 530 470 535
rect 425 495 440 530
rect 460 495 470 530
rect 425 490 470 495
rect 640 530 685 535
rect 640 495 650 530
rect 670 495 685 530
rect 640 490 685 495
rect 705 530 750 535
rect 705 495 720 530
rect 740 495 750 530
rect 705 490 750 495
rect 920 530 965 535
rect 920 495 930 530
rect 950 495 965 530
rect 920 490 965 495
rect 985 530 1030 535
rect 985 495 1000 530
rect 1020 495 1030 530
rect 985 490 1030 495
rect 1200 530 1245 535
rect 1200 495 1210 530
rect 1230 495 1245 530
rect 1200 490 1245 495
rect 1265 530 1310 535
rect 1265 495 1280 530
rect 1300 495 1310 530
rect 1265 490 1310 495
rect 1480 530 1525 535
rect 1480 495 1490 530
rect 1510 495 1525 530
rect 1480 490 1525 495
rect 1545 530 1590 535
rect 1545 495 1560 530
rect 1580 495 1590 530
rect 1545 490 1590 495
<< ndiffc >>
rect 90 385 110 420
rect 160 385 180 420
rect 370 385 390 420
rect 440 385 460 420
rect 650 385 670 420
rect 720 385 740 420
rect 930 385 950 420
rect 1000 385 1020 420
rect 1210 385 1230 420
rect 1280 385 1300 420
rect 1490 385 1510 420
rect 1560 385 1580 420
<< pdiffc >>
rect 90 495 110 530
rect 160 495 180 530
rect 370 495 390 530
rect 440 495 460 530
rect 650 495 670 530
rect 720 495 740 530
rect 930 495 950 530
rect 1000 495 1020 530
rect 1210 495 1230 530
rect 1280 495 1300 530
rect 1490 495 1510 530
rect 1560 495 1580 530
<< psubdiff >>
rect 80 315 95 345
rect 120 315 135 345
rect 360 315 375 345
rect 455 315 470 345
rect 640 315 655 345
rect 680 315 695 345
rect 920 315 935 345
rect 1015 315 1030 345
rect 1200 315 1215 345
rect 1240 315 1255 345
rect 1480 315 1495 345
rect 1575 315 1590 345
<< nsubdiff >>
rect 80 570 95 600
rect 120 570 135 600
rect 360 570 375 600
rect 455 570 470 600
rect 640 570 655 600
rect 680 570 695 600
rect 360 565 400 570
rect 920 570 935 600
rect 1015 570 1030 600
rect 1200 570 1215 600
rect 1240 570 1255 600
rect 920 565 960 570
rect 1480 570 1495 600
rect 1575 570 1590 600
rect 1480 565 1520 570
<< psubdiffcont >>
rect 95 315 120 345
rect 375 315 455 345
rect 655 315 680 345
rect 935 315 1015 345
rect 1215 315 1240 345
rect 1495 315 1575 345
<< nsubdiffcont >>
rect 95 570 120 600
rect 375 570 455 600
rect 655 570 680 600
rect 935 570 1015 600
rect 1215 570 1240 600
rect 1495 570 1575 600
<< poly >>
rect 155 595 210 600
rect 155 565 165 595
rect 200 565 210 595
rect 715 595 770 600
rect 715 565 725 595
rect 760 565 770 595
rect 1275 595 1330 600
rect 1275 565 1285 595
rect 1320 565 1330 595
rect 155 560 210 565
rect 715 560 770 565
rect 1275 560 1330 565
rect 125 545 210 560
rect 125 535 145 545
rect 405 535 425 550
rect 685 545 770 560
rect 685 535 705 545
rect 965 535 985 550
rect 1245 545 1330 560
rect 1245 535 1265 545
rect 1525 535 1545 550
rect 125 475 145 490
rect 405 475 425 490
rect 685 475 705 490
rect 965 475 985 490
rect 1245 475 1265 490
rect 1525 475 1545 490
rect 170 465 210 475
rect 170 445 175 465
rect 205 445 210 465
rect 125 425 145 440
rect 170 435 210 445
rect 340 465 425 475
rect 340 445 350 465
rect 395 445 425 465
rect 340 435 425 445
rect 730 465 770 475
rect 730 445 735 465
rect 765 445 770 465
rect 405 425 425 435
rect 685 425 705 440
rect 730 435 770 445
rect 900 465 985 475
rect 900 445 910 465
rect 955 445 985 465
rect 900 435 985 445
rect 1290 465 1330 475
rect 1290 445 1295 465
rect 1325 445 1330 465
rect 965 425 985 435
rect 1245 425 1265 440
rect 1290 435 1330 445
rect 1460 465 1545 475
rect 1460 445 1470 465
rect 1515 445 1545 465
rect 1460 435 1545 445
rect 1525 425 1545 435
rect 125 370 145 380
rect 125 355 210 370
rect 405 365 425 380
rect 685 370 705 380
rect 685 355 770 370
rect 965 365 985 380
rect 1245 370 1265 380
rect 1245 355 1330 370
rect 1525 365 1545 380
rect 155 350 210 355
rect 155 320 165 350
rect 200 320 210 350
rect 715 350 770 355
rect 155 315 210 320
rect 715 320 725 350
rect 760 320 770 350
rect 1275 350 1330 355
rect 715 315 770 320
rect 1275 320 1285 350
rect 1320 320 1330 350
rect 1275 315 1330 320
<< polycont >>
rect 165 565 200 595
rect 725 565 760 595
rect 1285 565 1320 595
rect 175 445 205 465
rect 350 445 395 465
rect 735 445 765 465
rect 910 445 955 465
rect 1295 445 1325 465
rect 1470 445 1515 465
rect 165 320 200 350
rect 725 320 760 350
rect 1285 320 1320 350
<< locali >>
rect 155 645 210 655
rect 155 625 160 645
rect 205 625 210 645
rect 80 595 95 600
rect 120 595 135 600
rect 80 575 90 595
rect 125 575 135 595
rect 80 570 95 575
rect 120 570 135 575
rect 155 595 210 625
rect 715 645 770 655
rect 715 625 720 645
rect 765 625 770 645
rect 155 565 165 595
rect 200 565 210 595
rect 155 560 210 565
rect 360 595 375 600
rect 455 595 470 600
rect 360 575 370 595
rect 460 575 470 595
rect 360 570 375 575
rect 455 570 470 575
rect 640 595 655 600
rect 680 595 695 600
rect 640 575 650 595
rect 685 575 695 595
rect 640 570 655 575
rect 680 570 695 575
rect 715 595 770 625
rect 1275 645 1330 655
rect 1275 625 1280 645
rect 1325 625 1330 645
rect 80 530 120 545
rect 80 495 90 530
rect 110 495 120 530
rect 80 475 120 495
rect 80 440 85 475
rect 115 440 120 475
rect 80 420 120 440
rect 80 385 90 420
rect 110 385 120 420
rect 80 380 120 385
rect 150 530 190 535
rect 150 495 160 530
rect 180 495 190 530
rect 150 475 190 495
rect 360 530 400 570
rect 640 560 680 570
rect 715 565 725 595
rect 760 565 770 595
rect 715 560 770 565
rect 920 595 935 600
rect 1015 595 1030 600
rect 920 575 930 595
rect 1020 575 1030 595
rect 920 570 935 575
rect 1015 570 1030 575
rect 1200 595 1215 600
rect 1240 595 1255 600
rect 1200 575 1210 595
rect 1245 575 1255 595
rect 1200 570 1215 575
rect 1240 570 1255 575
rect 1275 595 1330 625
rect 360 495 370 530
rect 390 495 400 530
rect 360 490 400 495
rect 430 530 470 535
rect 430 495 440 530
rect 460 495 470 530
rect 430 475 470 495
rect 150 440 160 475
rect 200 465 210 475
rect 205 445 210 465
rect 340 445 350 470
rect 395 445 405 470
rect 200 440 210 445
rect 150 435 210 440
rect 430 440 440 475
rect 150 420 190 435
rect 150 385 160 420
rect 180 385 190 420
rect 150 380 190 385
rect 360 420 400 425
rect 360 385 370 420
rect 390 385 400 420
rect 155 350 210 355
rect 80 340 95 345
rect 120 340 135 345
rect 80 320 90 340
rect 125 320 135 340
rect 80 315 95 320
rect 120 315 135 320
rect 155 320 165 350
rect 200 320 210 350
rect 155 295 210 320
rect 360 345 400 385
rect 430 420 470 440
rect 430 385 440 420
rect 460 385 470 420
rect 430 380 470 385
rect 640 530 680 535
rect 640 495 650 530
rect 670 495 680 530
rect 640 470 680 495
rect 675 445 680 470
rect 640 420 680 445
rect 640 385 650 420
rect 670 385 680 420
rect 640 380 680 385
rect 710 530 750 535
rect 710 495 720 530
rect 740 495 750 530
rect 710 475 750 495
rect 920 530 960 570
rect 1200 560 1240 570
rect 1275 565 1285 595
rect 1320 565 1330 595
rect 1275 560 1330 565
rect 1480 595 1495 600
rect 1575 595 1590 600
rect 1480 575 1490 595
rect 1580 575 1590 595
rect 1480 570 1495 575
rect 1575 570 1590 575
rect 920 495 930 530
rect 950 495 960 530
rect 920 490 960 495
rect 990 530 1030 535
rect 990 495 1000 530
rect 1020 495 1030 530
rect 990 475 1030 495
rect 710 470 770 475
rect 710 440 720 470
rect 760 465 770 470
rect 765 445 770 465
rect 900 445 910 470
rect 955 445 965 470
rect 760 440 770 445
rect 710 435 770 440
rect 990 440 1000 475
rect 710 420 750 435
rect 710 385 720 420
rect 740 385 750 420
rect 710 380 750 385
rect 920 420 960 425
rect 920 385 930 420
rect 950 385 960 420
rect 715 350 770 355
rect 360 340 375 345
rect 455 340 470 345
rect 360 320 370 340
rect 460 320 470 340
rect 360 315 375 320
rect 455 315 470 320
rect 640 340 655 345
rect 680 340 695 345
rect 640 320 650 340
rect 685 320 695 340
rect 640 315 655 320
rect 680 315 695 320
rect 715 320 725 350
rect 760 320 770 350
rect 155 265 165 295
rect 200 265 210 295
rect 155 260 210 265
rect 715 295 770 320
rect 920 345 960 385
rect 990 420 1030 440
rect 990 385 1000 420
rect 1020 385 1030 420
rect 990 380 1030 385
rect 1200 530 1240 535
rect 1200 495 1210 530
rect 1230 495 1240 530
rect 1200 470 1240 495
rect 1235 445 1240 470
rect 1200 420 1240 445
rect 1200 385 1210 420
rect 1230 385 1240 420
rect 1200 380 1240 385
rect 1270 530 1310 535
rect 1270 495 1280 530
rect 1300 495 1310 530
rect 1270 475 1310 495
rect 1480 530 1520 570
rect 1480 495 1490 530
rect 1510 495 1520 530
rect 1480 490 1520 495
rect 1550 530 1590 535
rect 1550 495 1560 530
rect 1580 495 1590 530
rect 1550 475 1590 495
rect 1270 470 1330 475
rect 1270 440 1280 470
rect 1320 465 1330 470
rect 1325 445 1330 465
rect 1460 445 1470 470
rect 1515 445 1525 470
rect 1320 440 1330 445
rect 1270 435 1330 440
rect 1550 440 1555 475
rect 1585 440 1590 475
rect 1270 420 1310 435
rect 1270 385 1280 420
rect 1300 385 1310 420
rect 1270 380 1310 385
rect 1480 420 1520 425
rect 1480 385 1490 420
rect 1510 385 1520 420
rect 1275 350 1330 355
rect 920 340 935 345
rect 1015 340 1030 345
rect 920 320 930 340
rect 1020 320 1030 340
rect 920 315 935 320
rect 1015 315 1030 320
rect 1200 340 1215 345
rect 1240 340 1255 345
rect 1200 320 1210 340
rect 1245 320 1255 340
rect 1200 315 1215 320
rect 1240 315 1255 320
rect 1275 320 1285 350
rect 1320 320 1330 350
rect 715 265 725 295
rect 760 265 770 295
rect 715 260 770 265
rect 1275 295 1330 320
rect 1480 345 1520 385
rect 1550 420 1590 440
rect 1550 385 1560 420
rect 1580 385 1590 420
rect 1550 380 1590 385
rect 1480 340 1495 345
rect 1575 340 1590 345
rect 1480 320 1490 340
rect 1580 320 1590 340
rect 1480 315 1495 320
rect 1575 315 1590 320
rect 1275 265 1285 295
rect 1320 265 1330 295
rect 1275 260 1330 265
<< viali >>
rect 160 625 205 645
rect 90 575 95 595
rect 95 575 120 595
rect 120 575 125 595
rect 720 625 765 645
rect 370 575 375 595
rect 375 575 455 595
rect 455 575 460 595
rect 650 575 655 595
rect 655 575 680 595
rect 680 575 685 595
rect 1280 625 1325 645
rect 85 440 115 475
rect 930 575 935 595
rect 935 575 1015 595
rect 1015 575 1020 595
rect 1210 575 1215 595
rect 1215 575 1240 595
rect 1240 575 1245 595
rect 160 465 200 475
rect 160 445 175 465
rect 175 445 200 465
rect 350 465 395 470
rect 350 445 395 465
rect 160 440 200 445
rect 440 440 470 475
rect 90 320 95 340
rect 95 320 120 340
rect 120 320 125 340
rect 640 445 675 470
rect 1490 575 1495 595
rect 1495 575 1575 595
rect 1575 575 1580 595
rect 720 465 760 470
rect 720 445 735 465
rect 735 445 760 465
rect 910 465 955 470
rect 910 445 955 465
rect 720 440 760 445
rect 1000 440 1030 475
rect 370 320 375 340
rect 375 320 455 340
rect 455 320 460 340
rect 650 320 655 340
rect 655 320 680 340
rect 680 320 685 340
rect 165 265 200 295
rect 1200 445 1235 470
rect 1280 465 1320 470
rect 1280 445 1295 465
rect 1295 445 1320 465
rect 1470 465 1515 470
rect 1470 445 1515 465
rect 1280 440 1320 445
rect 1555 440 1585 475
rect 930 320 935 340
rect 935 320 1015 340
rect 1015 320 1020 340
rect 1210 320 1215 340
rect 1215 320 1240 340
rect 1240 320 1245 340
rect 725 265 760 295
rect 1490 320 1495 340
rect 1495 320 1575 340
rect 1575 320 1580 340
rect 1285 265 1320 295
<< metal1 >>
rect 80 645 1330 655
rect 80 625 160 645
rect 205 625 720 645
rect 765 625 1280 645
rect 1325 625 1330 645
rect 80 615 1330 625
rect 80 595 1590 600
rect 80 575 90 595
rect 125 575 370 595
rect 460 575 650 595
rect 685 575 930 595
rect 1020 575 1210 595
rect 1245 575 1490 595
rect 1580 575 1590 595
rect 80 560 1590 575
rect 80 495 1590 535
rect 80 475 120 495
rect 1550 480 1590 495
rect 80 440 85 475
rect 115 440 120 475
rect 80 420 120 440
rect 150 475 210 480
rect 150 440 160 475
rect 200 440 210 475
rect 150 435 210 440
rect 340 470 405 480
rect 340 445 350 470
rect 395 445 405 470
rect 340 435 405 445
rect 430 475 680 480
rect 430 440 440 475
rect 470 470 680 475
rect 470 445 640 470
rect 675 445 680 470
rect 470 440 680 445
rect 430 435 680 440
rect 710 470 770 480
rect 710 440 720 470
rect 760 440 770 470
rect 710 435 770 440
rect 900 470 965 480
rect 900 445 910 470
rect 955 445 965 470
rect 900 435 965 445
rect 990 475 1240 480
rect 990 440 1000 475
rect 1030 470 1240 475
rect 1030 445 1200 470
rect 1235 445 1240 470
rect 1030 440 1240 445
rect 990 435 1240 440
rect 1270 470 1330 480
rect 1270 440 1280 470
rect 1320 440 1330 470
rect 1270 435 1330 440
rect 1460 470 1525 480
rect 1460 445 1470 470
rect 1515 445 1525 470
rect 1460 435 1525 445
rect 1550 475 1690 480
rect 1550 440 1555 475
rect 1585 440 1690 475
rect 1550 430 1690 440
rect 1550 420 1590 430
rect 80 380 1590 420
rect 80 340 1590 355
rect 80 320 90 340
rect 125 320 370 340
rect 460 320 650 340
rect 685 320 930 340
rect 1020 320 1210 340
rect 1245 320 1490 340
rect 1580 320 1590 340
rect 80 315 1590 320
rect 155 295 1330 300
rect 155 265 165 295
rect 200 265 725 295
rect 760 265 1285 295
rect 1320 265 1330 295
rect 155 260 1330 265
rect 1350 155 1590 315
rect 1350 -335 1360 155
rect 1580 -335 1590 155
rect 1350 -345 1590 -335
<< via1 >>
rect 210 435 340 480
rect 770 435 900 480
rect 1330 435 1460 480
rect 1360 -335 1580 155
<< metal2 >>
rect 200 435 210 480
rect 340 435 350 480
rect 760 435 770 480
rect 900 435 910 480
rect 1320 435 1330 480
rect 1460 435 1470 480
rect 1350 155 1590 165
rect 1350 -335 1360 155
rect 1580 -335 1590 155
rect 1350 -345 1590 -335
<< via2 >>
rect 210 440 340 480
rect 770 435 900 475
rect 1330 440 1460 480
rect 1360 -335 1580 155
<< metal3 >>
rect -300 725 745 1770
rect 905 730 1950 1775
rect 200 480 350 725
rect 1320 480 1470 730
rect 200 440 210 480
rect 340 440 350 480
rect 200 435 350 440
rect 760 475 910 480
rect 760 435 770 475
rect 900 435 910 475
rect 1320 440 1330 480
rect 1460 440 1470 480
rect 1320 435 1470 440
rect 760 185 910 435
rect 240 -855 1280 185
rect 1350 155 1590 165
rect 1350 -335 1360 155
rect 1580 -335 1590 155
rect 1350 -345 1590 -335
<< via3 >>
rect 1360 -335 1580 155
<< mimcap >>
rect -275 1210 725 1745
rect -275 760 -265 1210
rect 210 760 725 1210
rect -275 745 725 760
rect 925 1210 1925 1750
rect 925 760 935 1210
rect 1485 760 1925 1210
rect 925 750 1925 760
rect 260 150 1260 165
rect 260 -345 745 150
rect 1245 -345 1260 150
rect 260 -835 1260 -345
<< mimcapcontact >>
rect -265 760 210 1210
rect 935 760 1485 1210
rect 745 -345 1245 150
<< metal4 >>
rect -265 1210 210 1215
rect 210 760 935 1210
rect 1485 760 1925 1210
rect -265 755 210 760
rect 745 165 1245 760
rect 740 155 1590 165
rect 740 150 1360 155
rect 740 -345 745 150
rect 1245 -335 1360 150
rect 1580 -335 1590 155
rect 1245 -345 1590 -335
rect 740 -350 1260 -345
<< labels >>
flabel metal1 s 1590 581 1590 581 3 FreeSans 160 0 0 0 VPWR
port 0 e
flabel metal1 s 80 631 80 631 7 FreeSans 160 0 0 0 VCON-
port 1 w
flabel metal1 s 1690 454 1690 454 3 FreeSans 160 0 0 0 OUT_VCO
port 2 e
flabel metal1 s 156 277 156 277 7 FreeSans 160 0 0 0 VCON+
port 3 w
flabel metal1 s 1590 249 1590 249 3 FreeSans 160 0 0 0 VGND
port 4 e
<< end >>
