magic
tech sky130A
magscale 1 2
timestamp 1717247908
<< nwell >>
rect 580 238 3148 428
rect 582 -26 3148 238
<< pwell >>
rect 582 -498 3148 -88
rect 2152 -564 2224 -498
rect 2550 -502 2584 -498
<< pmos >>
rect 1636 40 1666 130
<< pdiff >>
rect 1578 40 1636 130
rect 1666 40 1724 130
<< psubdiff >>
rect 1230 -334 1288 -310
rect 1230 -400 1242 -334
rect 1276 -400 1288 -334
rect 1230 -424 1288 -400
rect 2450 -334 2508 -310
rect 2450 -400 2462 -334
rect 2496 -400 2508 -334
rect 2450 -424 2508 -400
<< nsubdiff >>
rect 1230 286 1288 310
rect 1230 220 1242 286
rect 1276 220 1288 286
rect 2450 286 2508 310
rect 1230 196 1288 220
rect 2450 220 2462 286
rect 2496 220 2508 286
rect 2450 196 2508 220
<< psubdiffcont >>
rect 1242 -400 1276 -334
rect 2462 -400 2496 -334
<< nsubdiffcont >>
rect 1242 220 1276 286
rect 2462 220 2496 286
<< poly >>
rect 1854 214 1922 224
rect 1854 178 1872 214
rect 1906 178 1922 214
rect 1854 156 1922 178
rect 602 74 636 114
rect 1200 -10 1230 156
rect 1636 130 1666 156
rect 1144 -26 1230 -10
rect 1636 -22 1666 40
rect 1854 14 1884 156
rect 1144 -60 1154 -26
rect 1190 -60 1230 -26
rect 1144 -76 1230 -60
rect 848 -134 918 -118
rect 848 -168 864 -134
rect 900 -168 918 -134
rect 848 -184 918 -168
rect 1200 -240 1230 -76
rect 1526 -38 1666 -22
rect 1526 -72 1542 -38
rect 1578 -56 1666 -38
rect 2290 -10 2320 156
rect 2508 -10 2538 156
rect 3092 54 3128 100
rect 2290 -26 2376 -10
rect 1578 -72 1594 -56
rect 1526 -88 1594 -72
rect 2290 -60 2326 -26
rect 2364 -60 2376 -26
rect 2290 -76 2376 -60
rect 2508 -26 2594 -10
rect 2508 -60 2544 -26
rect 2580 -60 2594 -26
rect 2508 -76 2594 -60
rect 2290 -240 2320 -76
rect 2508 -240 2538 -76
rect 2808 -132 2876 -116
rect 2808 -152 2824 -132
rect 2786 -166 2824 -152
rect 2860 -166 2876 -132
rect 2786 -182 2876 -166
rect 848 -256 1060 -240
rect 848 -290 864 -256
rect 900 -270 1060 -256
rect 1636 -256 1704 -240
rect 900 -290 916 -270
rect 848 -306 916 -290
rect 1636 -292 1652 -256
rect 1688 -292 1704 -256
rect 1636 -306 1704 -292
rect 1854 -256 1922 -240
rect 1854 -292 1870 -256
rect 1906 -292 1922 -256
rect 1854 -306 1922 -292
rect 2072 -256 2140 -240
rect 2072 -292 2088 -256
rect 2124 -292 2140 -256
rect 2072 -306 2140 -292
rect 2808 -256 2876 -240
rect 2808 -290 2824 -256
rect 2860 -290 2876 -256
rect 2808 -306 2876 -290
<< polycont >>
rect 1872 178 1906 214
rect 1154 -60 1190 -26
rect 864 -168 900 -134
rect 1542 -72 1578 -38
rect 2326 -60 2364 -26
rect 2544 -60 2580 -26
rect 2824 -166 2860 -132
rect 864 -290 900 -256
rect 1652 -292 1688 -256
rect 1870 -292 1906 -256
rect 2088 -292 2124 -256
rect 2824 -290 2860 -256
<< locali >>
rect 694 374 760 388
rect 694 340 708 374
rect 744 340 760 374
rect 600 -32 636 114
rect 694 108 760 340
rect 956 374 1022 388
rect 956 340 972 374
rect 1008 340 1022 374
rect 956 110 1022 340
rect 1138 374 1204 388
rect 1138 340 1154 374
rect 1190 340 1204 374
rect 1138 246 1204 340
rect 1242 374 1276 388
rect 1242 286 1276 340
rect 2462 374 2496 388
rect 1154 36 1188 246
rect 1242 196 1276 220
rect 1416 294 2104 328
rect 1416 178 1450 294
rect 1854 214 1922 224
rect 1854 178 1872 214
rect 1906 178 1922 214
rect 1854 176 1922 178
rect 2070 176 2104 294
rect 2462 286 2496 340
rect 2532 374 2598 388
rect 2532 340 2548 374
rect 2584 340 2598 374
rect 2532 246 2598 340
rect 2704 374 2770 388
rect 2704 340 2718 374
rect 2754 340 2770 374
rect 2462 196 2496 220
rect 1144 -26 1200 -10
rect 600 -68 900 -32
rect 864 -134 900 -68
rect 1144 -60 1154 -26
rect 1190 -60 1200 -26
rect 1144 -76 1200 -60
rect 610 -464 644 -134
rect 864 -184 900 -168
rect 1242 -204 1276 116
rect 1372 -26 1406 134
rect 1372 -218 1406 -60
rect 1460 -22 1494 134
rect 1590 118 1624 134
rect 1460 -38 1578 -22
rect 1460 -72 1542 -38
rect 1460 -88 1578 -72
rect 1678 -26 1712 134
rect 1460 -218 1494 -88
rect 864 -256 900 -240
rect 864 -306 900 -292
rect 1242 -334 1276 -310
rect 1242 -424 1276 -400
rect 1416 -384 1450 -252
rect 1560 -328 1594 -122
rect 1678 -218 1712 -60
rect 1896 -26 1930 134
rect 1774 -218 1842 -120
rect 1896 -218 1930 -60
rect 2026 -136 2060 134
rect 2114 -26 2148 134
rect 1964 -218 2060 -136
rect 2114 -218 2148 -60
rect 1636 -292 1652 -256
rect 1688 -292 1704 -256
rect 1774 -328 1808 -218
rect 1964 -256 1998 -218
rect 1854 -292 1870 -256
rect 1906 -292 1998 -256
rect 2072 -292 2088 -256
rect 2124 -292 2140 -256
rect 1594 -362 1808 -328
rect 1416 -418 1430 -384
rect 2088 -396 2124 -292
rect 1464 -418 2124 -396
rect 1416 -430 2124 -418
rect 2244 -464 2278 134
rect 2332 34 2366 102
rect 2326 -26 2364 -10
rect 2326 -76 2364 -60
rect 2332 -328 2366 -120
rect 2462 -218 2496 134
rect 2550 36 2584 246
rect 2704 110 2770 340
rect 2968 374 3034 388
rect 2968 340 2984 374
rect 3020 340 3034 374
rect 2968 110 3034 340
rect 2538 -24 2594 -10
rect 3092 -20 3128 116
rect 2538 -26 2546 -24
rect 2538 -60 2544 -26
rect 2582 -58 2594 -24
rect 2580 -60 2594 -58
rect 2538 -76 2594 -60
rect 2824 -56 3128 -20
rect 2462 -334 2496 -310
rect 2550 -328 2584 -120
rect 2824 -132 2860 -56
rect 2824 -182 2860 -166
rect 2824 -256 2860 -240
rect 2824 -306 2860 -290
rect 2462 -424 2496 -400
rect 3084 -464 3118 -134
rect 610 -498 3118 -464
<< viali >>
rect 708 340 744 374
rect 972 340 1008 374
rect 1154 340 1190 374
rect 1242 340 1276 374
rect 2462 340 2496 374
rect 1872 178 1906 212
rect 2548 340 2584 374
rect 2718 340 2754 374
rect 1154 -60 1190 -26
rect 1370 -60 1406 -26
rect 1678 -60 1712 -26
rect 864 -290 900 -256
rect 864 -292 900 -290
rect 1242 -400 1276 -334
rect 1896 -60 1930 -26
rect 2112 -60 2150 -26
rect 1652 -292 1688 -256
rect 1560 -362 1594 -328
rect 1430 -418 1464 -384
rect 2326 -60 2364 -26
rect 2984 340 3020 374
rect 2546 -26 2582 -24
rect 2546 -58 2580 -26
rect 2580 -58 2582 -26
rect 2332 -362 2366 -328
rect 2462 -400 2496 -334
rect 2824 -290 2860 -256
rect 2550 -362 2584 -328
<< metal1 >>
rect 370 388 570 528
rect 370 374 1300 388
rect 370 340 708 374
rect 744 340 972 374
rect 1008 340 1154 374
rect 1190 340 1242 374
rect 1276 340 1300 374
rect 370 328 1300 340
rect 1360 328 1732 388
rect 1792 374 3142 388
rect 1792 340 2462 374
rect 2496 340 2548 374
rect 2584 340 2718 374
rect 2754 340 2984 374
rect 3020 340 3142 374
rect 1792 328 3142 340
rect 1242 260 2366 294
rect 370 116 570 182
rect 1242 116 1276 260
rect 1726 226 1798 232
rect 1726 218 1732 226
rect 1400 164 1466 218
rect 1584 166 1732 218
rect 1792 166 1798 226
rect 370 50 652 116
rect 370 -18 570 50
rect 694 -106 760 56
rect 828 50 912 116
rect 828 -106 864 50
rect 594 -200 654 -134
rect 682 -140 864 -106
rect 956 -26 1022 56
rect 1584 40 1630 166
rect 1758 130 1798 166
rect 1854 212 1922 260
rect 2154 226 2226 232
rect 1854 178 1872 212
rect 1906 178 1922 212
rect 1854 164 1922 178
rect 2054 212 2120 218
rect 2154 212 2160 226
rect 2054 176 2160 212
rect 2054 164 2120 176
rect 2154 166 2160 176
rect 2220 166 2226 226
rect 2154 160 2226 166
rect 1758 40 1848 130
rect 2332 102 2366 260
rect 3152 116 3352 182
rect 1148 -26 1196 -10
rect 1364 -26 1412 -10
rect 1708 -12 1780 -6
rect 1708 -20 1714 -12
rect 956 -60 1154 -26
rect 1190 -60 1370 -26
rect 1406 -60 1412 -26
rect 956 -140 1022 -60
rect 1148 -76 1196 -60
rect 1364 -76 1412 -60
rect 1666 -26 1714 -20
rect 1666 -60 1678 -26
rect 1712 -60 1714 -26
rect 1666 -66 1714 -60
rect 1708 -72 1714 -66
rect 1774 -72 1780 -12
rect 1708 -78 1780 -72
rect 1828 -12 1936 -6
rect 1828 -72 1834 -12
rect 1894 -26 1936 -12
rect 2314 -18 2370 -14
rect 2538 -18 2590 -12
rect 2704 -18 2770 56
rect 2824 50 2894 116
rect 1894 -60 1896 -26
rect 1930 -60 1936 -26
rect 1894 -72 1936 -60
rect 2100 -24 2770 -18
rect 2100 -26 2546 -24
rect 2100 -60 2112 -26
rect 2150 -60 2326 -26
rect 2364 -58 2546 -26
rect 2582 -58 2770 -24
rect 2364 -60 2770 -58
rect 2100 -64 2770 -60
rect 2100 -66 2370 -64
rect 2314 -72 2370 -66
rect 2538 -70 2590 -64
rect 1828 -78 1936 -72
rect 682 -498 770 -190
rect 828 -240 864 -140
rect 828 -256 916 -240
rect 828 -292 864 -256
rect 900 -292 916 -256
rect 828 -306 916 -292
rect 944 -498 1034 -276
rect 1148 -498 1194 -122
rect 1400 -308 1466 -242
rect 1636 -256 1704 -244
rect 2462 -256 2496 -124
rect 2704 -140 2770 -64
rect 2860 -106 2894 50
rect 2968 -106 3034 56
rect 3076 50 3352 116
rect 3152 -18 3352 50
rect 2860 -140 3034 -106
rect 2860 -240 2894 -140
rect 1636 -292 1652 -256
rect 1688 -292 2496 -256
rect 2818 -256 2894 -240
rect 1636 -306 1704 -292
rect 1230 -334 1288 -326
rect 1230 -400 1242 -334
rect 1276 -400 1288 -334
rect 1554 -328 1600 -316
rect 2550 -322 2584 -316
rect 2326 -328 2372 -322
rect 1554 -362 1560 -328
rect 1594 -362 1600 -328
rect 1230 -410 1288 -400
rect 1410 -370 1482 -364
rect 1554 -368 1600 -362
rect 2320 -362 2332 -328
rect 2366 -362 2378 -328
rect 2320 -364 2378 -362
rect 2450 -334 2508 -324
rect 2326 -368 2372 -364
rect 1242 -498 1276 -410
rect 1410 -430 1416 -370
rect 1476 -430 1482 -370
rect 1410 -436 1482 -430
rect 1560 -498 1594 -368
rect 2332 -498 2366 -368
rect 2450 -400 2462 -334
rect 2496 -400 2508 -334
rect 2544 -328 2590 -322
rect 2544 -362 2550 -328
rect 2584 -362 2590 -328
rect 2544 -368 2590 -362
rect 2450 -408 2508 -400
rect 2462 -498 2496 -408
rect 2550 -498 2584 -368
rect 2692 -498 2782 -276
rect 2818 -290 2824 -256
rect 2860 -290 2894 -256
rect 2818 -306 2894 -290
rect 2956 -498 3046 -188
rect 3074 -200 3134 -134
rect 370 -558 2158 -498
rect 2218 -558 3142 -498
rect 370 -698 570 -558
rect 1542 -600 1742 -594
rect 1542 -660 1676 -600
rect 1736 -660 1742 -600
rect 1542 -794 1742 -660
rect 1866 -602 2066 -596
rect 1866 -662 1872 -602
rect 1932 -662 2066 -602
rect 1866 -796 2066 -662
<< via1 >>
rect 1300 328 1360 388
rect 1732 328 1792 388
rect 1732 166 1792 226
rect 2160 166 2220 226
rect 1714 -72 1774 -12
rect 1834 -72 1894 -12
rect 1416 -384 1476 -370
rect 1416 -418 1430 -384
rect 1430 -418 1464 -384
rect 1464 -418 1476 -384
rect 1416 -430 1476 -418
rect 2158 -558 2218 -498
rect 1676 -660 1736 -600
rect 1872 -662 1932 -602
<< metal2 >>
rect 1294 388 1366 394
rect 1294 328 1300 388
rect 1360 328 1366 388
rect 1294 322 1366 328
rect 1726 388 1798 394
rect 1726 328 1732 388
rect 1792 328 1798 388
rect 1726 322 1798 328
rect 1314 -384 1348 322
rect 1746 232 1780 322
rect 1726 226 1798 232
rect 1726 166 1732 226
rect 1792 166 1798 226
rect 1726 160 1798 166
rect 2154 226 2226 232
rect 2154 166 2160 226
rect 2220 166 2226 226
rect 2154 160 2226 166
rect 1708 -12 1780 -6
rect 1708 -72 1714 -12
rect 1774 -72 1780 -12
rect 1708 -78 1780 -72
rect 1828 -12 1900 -6
rect 1828 -72 1834 -12
rect 1894 -72 1900 -12
rect 1828 -78 1900 -72
rect 1410 -370 1482 -364
rect 1410 -384 1416 -370
rect 1314 -418 1416 -384
rect 1410 -430 1416 -418
rect 1476 -430 1482 -370
rect 1410 -436 1482 -430
rect 1708 -594 1742 -78
rect 1670 -600 1742 -594
rect 1670 -660 1676 -600
rect 1736 -660 1742 -600
rect 1670 -666 1742 -660
rect 1866 -596 1900 -78
rect 2172 -492 2206 160
rect 2152 -498 2224 -492
rect 2152 -558 2158 -498
rect 2218 -558 2224 -498
rect 2152 -564 2224 -558
rect 1866 -602 1938 -596
rect 1866 -662 1872 -602
rect 1932 -662 1938 -602
rect 1866 -668 1938 -662
use sky130_fd_pr__nfet_01v8_9NP8AN  sky130_fd_pr__nfet_01v8_9NP8AN_0
timestamp 1717214842
transform 1 0 2087 0 1 -169
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_VZM9AN  sky130_fd_pr__nfet_01v8_VZM9AN_0
timestamp 1717214842
transform -1 0 1215 0 -1 -169
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_27PL9K  sky130_fd_pr__pfet_01v8_27PL9K_0
timestamp 1717214842
transform -1 0 1215 0 -1 85
box -109 -107 109 107
use sky130_fd_pr__pfet_01v8_27PL9Z  sky130_fd_pr__pfet_01v8_27PL9Z_0
timestamp 1717214842
transform 0 1 953 -1 0 83
box -109 -109 109 143
use sky130_fd_pr__pfet_01v8_27PL9Z  sky130_fd_pr__pfet_01v8_27PL9Z_1
timestamp 1717214842
transform 0 1 691 -1 0 83
box -109 -109 109 143
use sky130_fd_pr__pfet_01v8_52DJGB  sky130_fd_pr__pfet_01v8_52DJGB_0
timestamp 1717182109
transform 1 0 1651 0 1 85
box -109 -107 109 107
use sky130_fd_pr__pfet_01v8_MJZT9K  sky130_fd_pr__pfet_01v8_MJZT9K_0
timestamp 1717214842
transform 1 0 2087 0 1 121
box -109 -143 109 109
use sky130_fd_pr__nfet_01v8_9NESAN  XM2
timestamp 1717214842
transform 0 1 696 -1 0 -167
box -73 -102 73 102
use sky130_fd_pr__nfet_01v8_9NP8AN  XM5
timestamp 1717214842
transform 0 1 989 -1 0 -167
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_9NP8AN  XM6
timestamp 1717214842
transform 0 1 989 -1 0 -255
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_52DJGB  XM8
timestamp 1717182109
transform 1 0 2305 0 1 85
box -109 -107 109 107
use sky130_fd_pr__nfet_01v8_BH4Y4M  XM9
timestamp 1717182109
transform 1 0 2305 0 1 -169
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_52DJGB  XM10
timestamp 1717182109
transform 1 0 2523 0 1 85
box -109 -107 109 107
use sky130_fd_pr__nfet_01v8_BH4Y4M  XM11
timestamp 1717182109
transform 1 0 2523 0 1 -169
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_AWEQGB  XM12
timestamp 1717230866
transform 0 1 2773 -1 0 83
box -109 -143 109 109
use sky130_fd_pr__nfet_01v8_BH4Y4M  XM13
timestamp 1717182109
transform 0 1 2737 -1 0 -167
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_AWEQGB  XM14
timestamp 1717230866
transform 0 1 3037 -1 0 83
box -109 -143 109 109
use sky130_fd_pr__nfet_01v8_ZVHWZ3  XM15
timestamp 1717230866
transform 0 1 3032 -1 0 -167
box -73 -102 73 102
use sky130_fd_pr__nfet_01v8_BH4Y4M  XM16
timestamp 1717182109
transform 0 1 2737 -1 0 -255
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_27PL9K  XM17
timestamp 1717214842
transform 1 0 1869 0 1 85
box -109 -107 109 107
use sky130_fd_pr__nfet_01v8_9NP8AN  XM18
timestamp 1717214842
transform 1 0 1869 0 1 -169
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_MJZT9K  XM19
timestamp 1717214842
transform 1 0 1433 0 1 121
box -109 -143 109 109
use sky130_fd_pr__nfet_01v8_9N7ETN  XM20
timestamp 1717230866
transform -1 0 1433 0 -1 -200
box -73 -102 73 102
use sky130_fd_pr__nfet_01v8_BH4Y4M  XM45
timestamp 1717182109
transform 1 0 1651 0 1 -169
box -73 -71 73 71
<< labels >>
flabel metal1 s 370 -612 370 -612 7 FreeSans 320 0 0 0 VN
port 0 w
flabel metal1 s 2066 -698 2066 -698 3 FreeSans 320 0 0 0 VCn
port 1 e
flabel metal1 s 370 78 370 78 7 FreeSans 320 0 0 0 REF
port 2 w
flabel metal1 s 3352 82 3352 82 3 FreeSans 320 0 0 0 FEEDBACK
port 3 e
flabel metal1 s 370 440 370 440 7 FreeSans 320 0 0 0 VP
port 4 w
flabel metal1 s 1542 -698 1542 -698 7 FreeSans 320 0 0 0 VCp
port 5 w
<< end >>
